LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY voltage2distance_long IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      voltage        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      distance       :  OUT   STD_LOGIC_VECTOR(12 DOWNTO 0));  
END voltage2distance_long;

ARCHITECTURE behavior OF voltage2distance_long IS

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 3393 ),
( 3385 ),
( 3377 ),
( 3369 ),
( 3361 ),
( 3353 ),
( 3345 ),
( 3337 ),
( 3329 ),
( 3322 ),
( 3314 ),
( 3306 ),
( 3298 ),
( 3291 ),
( 3283 ),
( 3276 ),
( 3268 ),
( 3260 ),
( 3253 ),
( 3245 ),
( 3238 ),
( 3230 ),
( 3223 ),
( 3216 ),
( 3208 ),
( 3201 ),
( 3194 ),
( 3186 ),
( 3179 ),
( 3172 ),
( 3165 ),
( 3158 ),
( 3150 ),
( 3143 ),
( 3136 ),
( 3129 ),
( 3122 ),
( 3115 ),
( 3108 ),
( 3101 ),
( 3094 ),
( 3087 ),
( 3080 ),
( 3074 ),
( 3067 ),
( 3060 ),
( 3053 ),
( 3046 ),
( 3040 ),
( 3033 ),
( 3026 ),
( 3020 ),
( 3013 ),
( 3006 ),
( 3000 ),
( 2993 ),
( 2987 ),
( 2980 ),
( 2974 ),
( 2967 ),
( 2961 ),
( 2954 ),
( 2948 ),
( 2942 ),
( 2935 ),
( 2929 ),
( 2923 ),
( 2916 ),
( 2910 ),
( 2904 ),
( 2898 ),
( 2891 ),
( 2885 ),
( 2879 ),
( 2873 ),
( 2867 ),
( 2861 ),
( 2855 ),
( 2849 ),
( 2843 ),
( 2837 ),
( 2831 ),
( 2825 ),
( 2819 ),
( 2813 ),
( 2807 ),
( 2801 ),
( 2795 ),
( 2790 ),
( 2784 ),
( 2778 ),
( 2772 ),
( 2767 ),
( 2761 ),
( 2755 ),
( 2750 ),
( 2744 ),
( 2738 ),
( 2733 ),
( 2727 ),
( 2722 ),
( 2716 ),
( 2710 ),
( 2705 ),
( 2699 ),
( 2694 ),
( 2689 ),
( 2683 ),
( 2678 ),
( 2672 ),
( 2667 ),
( 2662 ),
( 2656 ),
( 2651 ),
( 2646 ),
( 2640 ),
( 2635 ),
( 2630 ),
( 2625 ),
( 2620 ),
( 2614 ),
( 2609 ),
( 2604 ),
( 2599 ),
( 2594 ),
( 2589 ),
( 2584 ),
( 2579 ),
( 2574 ),
( 2569 ),
( 2564 ),
( 2559 ),
( 2554 ),
( 2549 ),
( 2544 ),
( 2539 ),
( 2534 ),
( 2529 ),
( 2524 ),
( 2519 ),
( 2515 ),
( 2510 ),
( 2505 ),
( 2500 ),
( 2496 ),
( 2491 ),
( 2486 ),
( 2481 ),
( 2477 ),
( 2472 ),
( 2467 ),
( 2463 ),
( 2458 ),
( 2454 ),
( 2449 ),
( 2444 ),
( 2440 ),
( 2435 ),
( 2431 ),
( 2426 ),
( 2422 ),
( 2417 ),
( 2413 ),
( 2408 ),
( 2404 ),
( 2400 ),
( 2395 ),
( 2391 ),
( 2386 ),
( 2382 ),
( 2378 ),
( 2373 ),
( 2369 ),
( 2365 ),
( 2361 ),
( 2356 ),
( 2352 ),
( 2348 ),
( 2344 ),
( 2339 ),
( 2335 ),
( 2331 ),
( 2327 ),
( 2323 ),
( 2319 ),
( 2314 ),
( 2310 ),
( 2306 ),
( 2302 ),
( 2298 ),
( 2294 ),
( 2290 ),
( 2286 ),
( 2282 ),
( 2278 ),
( 2274 ),
( 2270 ),
( 2266 ),
( 2262 ),
( 2258 ),
( 2254 ),
( 2250 ),
( 2247 ),
( 2243 ),
( 2239 ),
( 2235 ),
( 2231 ),
( 2227 ),
( 2224 ),
( 2220 ),
( 2216 ),
( 2212 ),
( 2208 ),
( 2205 ),
( 2201 ),
( 2197 ),
( 2194 ),
( 2190 ),
( 2186 ),
( 2183 ),
( 2179 ),
( 2175 ),
( 2172 ),
( 2168 ),
( 2164 ),
( 2161 ),
( 2157 ),
( 2154 ),
( 2150 ),
( 2147 ),
( 2143 ),
( 2140 ),
( 2136 ),
( 2132 ),
( 2129 ),
( 2126 ),
( 2122 ),
( 2119 ),
( 2115 ),
( 2112 ),
( 2108 ),
( 2105 ),
( 2101 ),
( 2098 ),
( 2095 ),
( 2091 ),
( 2088 ),
( 2085 ),
( 2081 ),
( 2078 ),
( 2075 ),
( 2071 ),
( 2068 ),
( 2065 ),
( 2062 ),
( 2058 ),
( 2055 ),
( 2052 ),
( 2049 ),
( 2045 ),
( 2042 ),
( 2039 ),
( 2036 ),
( 2033 ),
( 2029 ),
( 2026 ),
( 2023 ),
( 2020 ),
( 2017 ),
( 2014 ),
( 2011 ),
( 2008 ),
( 2004 ),
( 2001 ),
( 1998 ),
( 1995 ),
( 1992 ),
( 1989 ),
( 1986 ),
( 1983 ),
( 1980 ),
( 1977 ),
( 1974 ),
( 1971 ),
( 1968 ),
( 1965 ),
( 1962 ),
( 1959 ),
( 1956 ),
( 1953 ),
( 1951 ),
( 1948 ),
( 1945 ),
( 1942 ),
( 1939 ),
( 1936 ),
( 1933 ),
( 1930 ),
( 1927 ),
( 1925 ),
( 1922 ),
( 1919 ),
( 1916 ),
( 1913 ),
( 1911 ),
( 1908 ),
( 1905 ),
( 1902 ),
( 1899 ),
( 1897 ),
( 1894 ),
( 1891 ),
( 1888 ),
( 1886 ),
( 1883 ),
( 1880 ),
( 1878 ),
( 1875 ),
( 1872 ),
( 1870 ),
( 1867 ),
( 1864 ),
( 1862 ),
( 1859 ),
( 1856 ),
( 1854 ),
( 1851 ),
( 1848 ),
( 1846 ),
( 1843 ),
( 1841 ),
( 1838 ),
( 1835 ),
( 1833 ),
( 1830 ),
( 1828 ),
( 1825 ),
( 1823 ),
( 1820 ),
( 1818 ),
( 1815 ),
( 1813 ),
( 1810 ),
( 1808 ),
( 1805 ),
( 1803 ),
( 1800 ),
( 1798 ),
( 1795 ),
( 1793 ),
( 1790 ),
( 1788 ),
( 1785 ),
( 1783 ),
( 1781 ),
( 1778 ),
( 1776 ),
( 1773 ),
( 1771 ),
( 1769 ),
( 1766 ),
( 1764 ),
( 1762 ),
( 1759 ),
( 1757 ),
( 1754 ),
( 1752 ),
( 1750 ),
( 1747 ),
( 1745 ),
( 1743 ),
( 1740 ),
( 1738 ),
( 1736 ),
( 1734 ),
( 1731 ),
( 1729 ),
( 1727 ),
( 1724 ),
( 1722 ),
( 1720 ),
( 1718 ),
( 1715 ),
( 1713 ),
( 1711 ),
( 1709 ),
( 1707 ),
( 1704 ),
( 1702 ),
( 1700 ),
( 1698 ),
( 1696 ),
( 1693 ),
( 1691 ),
( 1689 ),
( 1687 ),
( 1685 ),
( 1683 ),
( 1680 ),
( 1678 ),
( 1676 ),
( 1674 ),
( 1672 ),
( 1670 ),
( 1668 ),
( 1665 ),
( 1663 ),
( 1661 ),
( 1659 ),
( 1657 ),
( 1655 ),
( 1653 ),
( 1651 ),
( 1649 ),
( 1647 ),
( 1645 ),
( 1643 ),
( 1640 ),
( 1638 ),
( 1636 ),
( 1634 ),
( 1632 ),
( 1630 ),
( 1628 ),
( 1626 ),
( 1624 ),
( 1622 ),
( 1620 ),
( 1618 ),
( 1616 ),
( 1614 ),
( 1612 ),
( 1610 ),
( 1608 ),
( 1606 ),
( 1604 ),
( 1602 ),
( 1600 ),
( 1599 ),
( 1597 ),
( 1595 ),
( 1593 ),
( 1591 ),
( 1589 ),
( 1587 ),
( 1585 ),
( 1583 ),
( 1581 ),
( 1579 ),
( 1577 ),
( 1575 ),
( 1574 ),
( 1572 ),
( 1570 ),
( 1568 ),
( 1566 ),
( 1564 ),
( 1562 ),
( 1560 ),
( 1559 ),
( 1557 ),
( 1555 ),
( 1553 ),
( 1551 ),
( 1549 ),
( 1548 ),
( 1546 ),
( 1544 ),
( 1542 ),
( 1540 ),
( 1538 ),
( 1537 ),
( 1535 ),
( 1533 ),
( 1531 ),
( 1529 ),
( 1528 ),
( 1526 ),
( 1524 ),
( 1522 ),
( 1521 ),
( 1519 ),
( 1517 ),
( 1515 ),
( 1513 ),
( 1512 ),
( 1510 ),
( 1508 ),
( 1506 ),
( 1505 ),
( 1503 ),
( 1501 ),
( 1500 ),
( 1498 ),
( 1496 ),
( 1494 ),
( 1493 ),
( 1491 ),
( 1489 ),
( 1488 ),
( 1486 ),
( 1484 ),
( 1482 ),
( 1481 ),
( 1479 ),
( 1477 ),
( 1476 ),
( 1474 ),
( 1472 ),
( 1471 ),
( 1469 ),
( 1467 ),
( 1466 ),
( 1464 ),
( 1462 ),
( 1461 ),
( 1459 ),
( 1458 ),
( 1456 ),
( 1454 ),
( 1453 ),
( 1451 ),
( 1449 ),
( 1448 ),
( 1446 ),
( 1445 ),
( 1443 ),
( 1441 ),
( 1440 ),
( 1438 ),
( 1436 ),
( 1435 ),
( 1433 ),
( 1432 ),
( 1430 ),
( 1429 ),
( 1427 ),
( 1425 ),
( 1424 ),
( 1422 ),
( 1421 ),
( 1419 ),
( 1418 ),
( 1416 ),
( 1414 ),
( 1413 ),
( 1411 ),
( 1410 ),
( 1408 ),
( 1407 ),
( 1405 ),
( 1404 ),
( 1402 ),
( 1401 ),
( 1399 ),
( 1398 ),
( 1396 ),
( 1394 ),
( 1393 ),
( 1391 ),
( 1390 ),
( 1388 ),
( 1387 ),
( 1385 ),
( 1384 ),
( 1382 ),
( 1381 ),
( 1379 ),
( 1378 ),
( 1376 ),
( 1375 ),
( 1374 ),
( 1372 ),
( 1371 ),
( 1369 ),
( 1368 ),
( 1366 ),
( 1365 ),
( 1363 ),
( 1362 ),
( 1360 ),
( 1359 ),
( 1357 ),
( 1356 ),
( 1355 ),
( 1353 ),
( 1352 ),
( 1350 ),
( 1349 ),
( 1347 ),
( 1346 ),
( 1344 ),
( 1343 ),
( 1342 ),
( 1340 ),
( 1339 ),
( 1337 ),
( 1336 ),
( 1335 ),
( 1333 ),
( 1332 ),
( 1330 ),
( 1329 ),
( 1328 ),
( 1326 ),
( 1325 ),
( 1323 ),
( 1322 ),
( 1321 ),
( 1319 ),
( 1318 ),
( 1316 ),
( 1315 ),
( 1314 ),
( 1312 ),
( 1311 ),
( 1310 ),
( 1308 ),
( 1307 ),
( 1305 ),
( 1304 ),
( 1303 ),
( 1301 ),
( 1300 ),
( 1299 ),
( 1297 ),
( 1296 ),
( 1295 ),
( 1293 ),
( 1292 ),
( 1291 ),
( 1289 ),
( 1288 ),
( 1287 ),
( 1285 ),
( 1284 ),
( 1283 ),
( 1281 ),
( 1280 ),
( 1279 ),
( 1277 ),
( 1276 ),
( 1275 ),
( 1273 ),
( 1272 ),
( 1271 ),
( 1270 ),
( 1268 ),
( 1267 ),
( 1266 ),
( 1264 ),
( 1263 ),
( 1262 ),
( 1261 ),
( 1259 ),
( 1258 ),
( 1257 ),
( 1255 ),
( 1254 ),
( 1253 ),
( 1252 ),
( 1250 ),
( 1249 ),
( 1248 ),
( 1246 ),
( 1245 ),
( 1244 ),
( 1243 ),
( 1241 ),
( 1240 ),
( 1239 ),
( 1238 ),
( 1236 ),
( 1235 ),
( 1234 ),
( 1233 ),
( 1231 ),
( 1230 ),
( 1229 ),
( 1228 ),
( 1227 ),
( 1225 ),
( 1224 ),
( 1223 ),
( 1222 ),
( 1220 ),
( 1219 ),
( 1218 ),
( 1217 ),
( 1216 ),
( 1214 ),
( 1213 ),
( 1212 ),
( 1211 ),
( 1209 ),
( 1208 ),
( 1207 ),
( 1206 ),
( 1205 ),
( 1203 ),
( 1202 ),
( 1201 ),
( 1200 ),
( 1199 ),
( 1197 ),
( 1196 ),
( 1195 ),
( 1194 ),
( 1193 ),
( 1192 ),
( 1190 ),
( 1189 ),
( 1188 ),
( 1187 ),
( 1186 ),
( 1185 ),
( 1183 ),
( 1182 ),
( 1181 ),
( 1180 ),
( 1179 ),
( 1178 ),
( 1176 ),
( 1175 ),
( 1174 ),
( 1173 ),
( 1172 ),
( 1171 ),
( 1170 ),
( 1168 ),
( 1167 ),
( 1166 ),
( 1165 ),
( 1164 ),
( 1163 ),
( 1162 ),
( 1160 ),
( 1159 ),
( 1158 ),
( 1157 ),
( 1156 ),
( 1155 ),
( 1154 ),
( 1153 ),
( 1151 ),
( 1150 ),
( 1149 ),
( 1148 ),
( 1147 ),
( 1146 ),
( 1145 ),
( 1144 ),
( 1143 ),
( 1141 ),
( 1140 ),
( 1139 ),
( 1138 ),
( 1137 ),
( 1136 ),
( 1135 ),
( 1134 ),
( 1133 ),
( 1132 ),
( 1130 ),
( 1129 ),
( 1128 ),
( 1127 ),
( 1126 ),
( 1125 ),
( 1124 ),
( 1123 ),
( 1122 ),
( 1121 ),
( 1120 ),
( 1119 ),
( 1118 ),
( 1117 ),
( 1115 ),
( 1114 ),
( 1113 ),
( 1112 ),
( 1111 ),
( 1110 ),
( 1109 ),
( 1108 ),
( 1107 ),
( 1106 ),
( 1105 ),
( 1104 ),
( 1103 ),
( 1102 ),
( 1101 ),
( 1100 ),
( 1099 ),
( 1098 ),
( 1097 ),
( 1096 ),
( 1094 ),
( 1093 ),
( 1092 ),
( 1091 ),
( 1090 ),
( 1089 ),
( 1088 ),
( 1087 ),
( 1086 ),
( 1085 ),
( 1084 ),
( 1083 ),
( 1082 ),
( 1081 ),
( 1080 ),
( 1079 ),
( 1078 ),
( 1077 ),
( 1076 ),
( 1075 ),
( 1074 ),
( 1073 ),
( 1072 ),
( 1071 ),
( 1070 ),
( 1069 ),
( 1068 ),
( 1067 ),
( 1066 ),
( 1065 ),
( 1064 ),
( 1063 ),
( 1062 ),
( 1061 ),
( 1060 ),
( 1059 ),
( 1058 ),
( 1057 ),
( 1056 ),
( 1055 ),
( 1054 ),
( 1053 ),
( 1052 ),
( 1052 ),
( 1051 ),
( 1050 ),
( 1049 ),
( 1048 ),
( 1047 ),
( 1046 ),
( 1045 ),
( 1044 ),
( 1043 ),
( 1042 ),
( 1041 ),
( 1040 ),
( 1039 ),
( 1038 ),
( 1037 ),
( 1036 ),
( 1035 ),
( 1034 ),
( 1033 ),
( 1032 ),
( 1032 ),
( 1031 ),
( 1030 ),
( 1029 ),
( 1028 ),
( 1027 ),
( 1026 ),
( 1025 ),
( 1024 ),
( 1023 ),
( 1022 ),
( 1021 ),
( 1020 ),
( 1019 ),
( 1019 ),
( 1018 ),
( 1017 ),
( 1016 ),
( 1015 ),
( 1014 ),
( 1013 ),
( 1012 ),
( 1011 ),
( 1010 ),
( 1009 ),
( 1009 ),
( 1008 ),
( 1007 ),
( 1006 ),
( 1005 ),
( 1004 ),
( 1003 ),
( 1002 ),
( 1001 ),
( 1001 ),
( 1000 ),
( 999 ),
( 998 ),
( 997 ),
( 996 ),
( 995 ),
( 994 ),
( 993 ),
( 993 ),
( 992 ),
( 991 ),
( 990 ),
( 989 ),
( 988 ),
( 987 ),
( 986 ),
( 986 ),
( 985 ),
( 984 ),
( 983 ),
( 982 ),
( 981 ),
( 980 ),
( 980 ),
( 979 ),
( 978 ),
( 977 ),
( 976 ),
( 975 ),
( 974 ),
( 974 ),
( 973 ),
( 972 ),
( 971 ),
( 970 ),
( 969 ),
( 969 ),
( 968 ),
( 967 ),
( 966 ),
( 965 ),
( 964 ),
( 964 ),
( 963 ),
( 962 ),
( 961 ),
( 960 ),
( 959 ),
( 959 ),
( 958 ),
( 957 ),
( 956 ),
( 955 ),
( 955 ),
( 954 ),
( 953 ),
( 952 ),
( 951 ),
( 951 ),
( 950 ),
( 949 ),
( 948 ),
( 947 ),
( 946 ),
( 946 ),
( 945 ),
( 944 ),
( 943 ),
( 943 ),
( 942 ),
( 941 ),
( 940 ),
( 939 ),
( 939 ),
( 938 ),
( 937 ),
( 936 ),
( 935 ),
( 935 ),
( 934 ),
( 933 ),
( 932 ),
( 932 ),
( 931 ),
( 930 ),
( 929 ),
( 928 ),
( 928 ),
( 927 ),
( 926 ),
( 925 ),
( 925 ),
( 924 ),
( 923 ),
( 922 ),
( 922 ),
( 921 ),
( 920 ),
( 919 ),
( 919 ),
( 918 ),
( 917 ),
( 916 ),
( 916 ),
( 915 ),
( 914 ),
( 913 ),
( 913 ),
( 912 ),
( 911 ),
( 910 ),
( 910 ),
( 909 ),
( 908 ),
( 907 ),
( 907 ),
( 906 ),
( 905 ),
( 904 ),
( 904 ),
( 903 ),
( 902 ),
( 902 ),
( 901 ),
( 900 ),
( 899 ),
( 899 ),
( 898 ),
( 897 ),
( 896 ),
( 896 ),
( 895 ),
( 894 ),
( 894 ),
( 893 ),
( 892 ),
( 892 ),
( 891 ),
( 890 ),
( 889 ),
( 889 ),
( 888 ),
( 887 ),
( 887 ),
( 886 ),
( 885 ),
( 884 ),
( 884 ),
( 883 ),
( 882 ),
( 882 ),
( 881 ),
( 880 ),
( 880 ),
( 879 ),
( 878 ),
( 878 ),
( 877 ),
( 876 ),
( 876 ),
( 875 ),
( 874 ),
( 874 ),
( 873 ),
( 872 ),
( 872 ),
( 871 ),
( 870 ),
( 870 ),
( 869 ),
( 868 ),
( 868 ),
( 867 ),
( 866 ),
( 866 ),
( 865 ),
( 864 ),
( 864 ),
( 863 ),
( 862 ),
( 862 ),
( 861 ),
( 860 ),
( 860 ),
( 859 ),
( 858 ),
( 858 ),
( 857 ),
( 856 ),
( 856 ),
( 855 ),
( 854 ),
( 854 ),
( 853 ),
( 853 ),
( 852 ),
( 851 ),
( 851 ),
( 850 ),
( 849 ),
( 849 ),
( 848 ),
( 847 ),
( 847 ),
( 846 ),
( 846 ),
( 845 ),
( 844 ),
( 844 ),
( 843 ),
( 842 ),
( 842 ),
( 841 ),
( 841 ),
( 840 ),
( 839 ),
( 839 ),
( 838 ),
( 838 ),
( 837 ),
( 836 ),
( 836 ),
( 835 ),
( 835 ),
( 834 ),
( 833 ),
( 833 ),
( 832 ),
( 832 ),
( 831 ),
( 830 ),
( 830 ),
( 829 ),
( 829 ),
( 828 ),
( 827 ),
( 827 ),
( 826 ),
( 826 ),
( 825 ),
( 824 ),
( 824 ),
( 823 ),
( 823 ),
( 822 ),
( 822 ),
( 821 ),
( 820 ),
( 820 ),
( 819 ),
( 819 ),
( 818 ),
( 817 ),
( 817 ),
( 816 ),
( 816 ),
( 815 ),
( 815 ),
( 814 ),
( 813 ),
( 813 ),
( 812 ),
( 812 ),
( 811 ),
( 811 ),
( 810 ),
( 810 ),
( 809 ),
( 808 ),
( 808 ),
( 807 ),
( 807 ),
( 806 ),
( 806 ),
( 805 ),
( 805 ),
( 804 ),
( 803 ),
( 803 ),
( 802 ),
( 802 ),
( 801 ),
( 801 ),
( 800 ),
( 800 ),
( 799 ),
( 799 ),
( 798 ),
( 798 ),
( 797 ),
( 796 ),
( 796 ),
( 795 ),
( 795 ),
( 794 ),
( 794 ),
( 793 ),
( 793 ),
( 792 ),
( 792 ),
( 791 ),
( 791 ),
( 790 ),
( 790 ),
( 789 ),
( 789 ),
( 788 ),
( 788 ),
( 787 ),
( 786 ),
( 786 ),
( 785 ),
( 785 ),
( 784 ),
( 784 ),
( 783 ),
( 783 ),
( 782 ),
( 782 ),
( 781 ),
( 781 ),
( 780 ),
( 780 ),
( 779 ),
( 779 ),
( 778 ),
( 778 ),
( 777 ),
( 777 ),
( 776 ),
( 776 ),
( 775 ),
( 775 ),
( 774 ),
( 774 ),
( 773 ),
( 773 ),
( 772 ),
( 772 ),
( 771 ),
( 771 ),
( 770 ),
( 770 ),
( 769 ),
( 769 ),
( 768 ),
( 768 ),
( 768 ),
( 767 ),
( 767 ),
( 766 ),
( 766 ),
( 765 ),
( 765 ),
( 764 ),
( 764 ),
( 763 ),
( 763 ),
( 762 ),
( 762 ),
( 761 ),
( 761 ),
( 760 ),
( 760 ),
( 759 ),
( 759 ),
( 759 ),
( 758 ),
( 758 ),
( 757 ),
( 757 ),
( 756 ),
( 756 ),
( 755 ),
( 755 ),
( 754 ),
( 754 ),
( 753 ),
( 753 ),
( 753 ),
( 752 ),
( 752 ),
( 751 ),
( 751 ),
( 750 ),
( 750 ),
( 749 ),
( 749 ),
( 748 ),
( 748 ),
( 748 ),
( 747 ),
( 747 ),
( 746 ),
( 746 ),
( 745 ),
( 745 ),
( 744 ),
( 744 ),
( 744 ),
( 743 ),
( 743 ),
( 742 ),
( 742 ),
( 741 ),
( 741 ),
( 741 ),
( 740 ),
( 740 ),
( 739 ),
( 739 ),
( 738 ),
( 738 ),
( 737 ),
( 737 ),
( 737 ),
( 736 ),
( 736 ),
( 735 ),
( 735 ),
( 735 ),
( 734 ),
( 734 ),
( 733 ),
( 733 ),
( 732 ),
( 732 ),
( 732 ),
( 731 ),
( 731 ),
( 730 ),
( 730 ),
( 729 ),
( 729 ),
( 729 ),
( 728 ),
( 728 ),
( 727 ),
( 727 ),
( 727 ),
( 726 ),
( 726 ),
( 725 ),
( 725 ),
( 724 ),
( 724 ),
( 724 ),
( 723 ),
( 723 ),
( 722 ),
( 722 ),
( 722 ),
( 721 ),
( 721 ),
( 720 ),
( 720 ),
( 720 ),
( 719 ),
( 719 ),
( 718 ),
( 718 ),
( 718 ),
( 717 ),
( 717 ),
( 716 ),
( 716 ),
( 716 ),
( 715 ),
( 715 ),
( 714 ),
( 714 ),
( 714 ),
( 713 ),
( 713 ),
( 712 ),
( 712 ),
( 712 ),
( 711 ),
( 711 ),
( 710 ),
( 710 ),
( 710 ),
( 709 ),
( 709 ),
( 709 ),
( 708 ),
( 708 ),
( 707 ),
( 707 ),
( 707 ),
( 706 ),
( 706 ),
( 705 ),
( 705 ),
( 705 ),
( 704 ),
( 704 ),
( 704 ),
( 703 ),
( 703 ),
( 702 ),
( 702 ),
( 702 ),
( 701 ),
( 701 ),
( 701 ),
( 700 ),
( 700 ),
( 699 ),
( 699 ),
( 699 ),
( 698 ),
( 698 ),
( 698 ),
( 697 ),
( 697 ),
( 696 ),
( 696 ),
( 696 ),
( 695 ),
( 695 ),
( 695 ),
( 694 ),
( 694 ),
( 693 ),
( 693 ),
( 693 ),
( 692 ),
( 692 ),
( 692 ),
( 691 ),
( 691 ),
( 691 ),
( 690 ),
( 690 ),
( 689 ),
( 689 ),
( 689 ),
( 688 ),
( 688 ),
( 688 ),
( 687 ),
( 687 ),
( 687 ),
( 686 ),
( 686 ),
( 685 ),
( 685 ),
( 685 ),
( 684 ),
( 684 ),
( 684 ),
( 683 ),
( 683 ),
( 683 ),
( 682 ),
( 682 ),
( 682 ),
( 681 ),
( 681 ),
( 680 ),
( 680 ),
( 680 ),
( 679 ),
( 679 ),
( 679 ),
( 678 ),
( 678 ),
( 678 ),
( 677 ),
( 677 ),
( 677 ),
( 676 ),
( 676 ),
( 675 ),
( 675 ),
( 675 ),
( 674 ),
( 674 ),
( 674 ),
( 673 ),
( 673 ),
( 673 ),
( 672 ),
( 672 ),
( 672 ),
( 671 ),
( 671 ),
( 671 ),
( 670 ),
( 670 ),
( 670 ),
( 669 ),
( 669 ),
( 669 ),
( 668 ),
( 668 ),
( 668 ),
( 667 ),
( 667 ),
( 666 ),
( 666 ),
( 666 ),
( 665 ),
( 665 ),
( 665 ),
( 664 ),
( 664 ),
( 664 ),
( 663 ),
( 663 ),
( 663 ),
( 662 ),
( 662 ),
( 662 ),
( 661 ),
( 661 ),
( 661 ),
( 660 ),
( 660 ),
( 660 ),
( 659 ),
( 659 ),
( 659 ),
( 658 ),
( 658 ),
( 658 ),
( 657 ),
( 657 ),
( 657 ),
( 656 ),
( 656 ),
( 656 ),
( 655 ),
( 655 ),
( 655 ),
( 654 ),
( 654 ),
( 654 ),
( 653 ),
( 653 ),
( 653 ),
( 652 ),
( 652 ),
( 652 ),
( 651 ),
( 651 ),
( 651 ),
( 650 ),
( 650 ),
( 650 ),
( 649 ),
( 649 ),
( 649 ),
( 648 ),
( 648 ),
( 647 ),
( 647 ),
( 647 ),
( 646 ),
( 646 ),
( 646 ),
( 645 ),
( 645 ),
( 645 ),
( 644 ),
( 644 ),
( 644 ),
( 643 ),
( 643 ),
( 643 ),
( 642 ),
( 642 ),
( 642 ),
( 641 ),
( 641 ),
( 641 ),
( 641 ),
( 640 ),
( 640 ),
( 640 ),
( 639 ),
( 639 ),
( 639 ),
( 638 ),
( 638 ),
( 638 ),
( 637 ),
( 637 ),
( 637 ),
( 636 ),
( 636 ),
( 636 ),
( 635 ),
( 635 ),
( 635 ),
( 634 ),
( 634 ),
( 634 ),
( 633 ),
( 633 ),
( 633 ),
( 632 ),
( 632 ),
( 632 ),
( 631 ),
( 631 ),
( 631 ),
( 630 ),
( 630 ),
( 630 ),
( 629 ),
( 629 ),
( 629 ),
( 628 ),
( 628 ),
( 628 ),
( 627 ),
( 627 ),
( 627 ),
( 626 ),
( 626 ),
( 626 ),
( 625 ),
( 625 ),
( 625 ),
( 624 ),
( 624 ),
( 624 ),
( 623 ),
( 623 ),
( 623 ),
( 622 ),
( 622 ),
( 622 ),
( 621 ),
( 621 ),
( 621 ),
( 620 ),
( 620 ),
( 620 ),
( 619 ),
( 619 ),
( 619 ),
( 618 ),
( 618 ),
( 618 ),
( 617 ),
( 617 ),
( 617 ),
( 616 ),
( 616 ),
( 616 ),
( 615 ),
( 615 ),
( 615 ),
( 614 ),
( 614 ),
( 614 ),
( 613 ),
( 613 ),
( 613 ),
( 612 ),
( 612 ),
( 612 ),
( 611 ),
( 611 ),
( 611 ),
( 610 ),
( 610 ),
( 610 ),
( 609 ),
( 609 ),
( 609 ),
( 608 ),
( 608 ),
( 608 ),
( 607 ),
( 607 ),
( 607 ),
( 606 ),
( 606 ),
( 606 ),
( 605 ),
( 605 ),
( 605 ),
( 604 ),
( 604 ),
( 604 ),
( 603 ),
( 603 ),
( 603 ),
( 602 ),
( 602 ),
( 602 ),
( 601 ),
( 601 ),
( 601 ),
( 600 ),
( 600 ),
( 600 ),
( 599 ),
( 599 ),
( 599 ),
( 598 ),
( 598 ),
( 598 ),
( 597 ),
( 597 ),
( 597 ),
( 596 ),
( 596 ),
( 596 ),
( 595 ),
( 595 ),
( 595 ),
( 594 ),
( 594 ),
( 594 ),
( 593 ),
( 593 ),
( 593 ),
( 592 ),
( 592 ),
( 592 ),
( 591 ),
( 591 ),
( 591 ),
( 590 ),
( 590 ),
( 590 ),
( 589 ),
( 589 ),
( 589 ),
( 588 ),
( 588 ),
( 588 ),
( 587 ),
( 587 ),
( 587 ),
( 586 ),
( 586 ),
( 586 ),
( 585 ),
( 585 ),
( 585 ),
( 584 ),
( 584 ),
( 584 ),
( 583 ),
( 583 ),
( 583 ),
( 582 ),
( 582 ),
( 582 ),
( 581 ),
( 581 ),
( 581 ),
( 580 ),
( 580 ),
( 580 ),
( 579 ),
( 579 ),
( 579 ),
( 578 ),
( 578 ),
( 578 ),
( 577 ),
( 577 ),
( 577 ),
( 576 ),
( 576 ),
( 576 ),
( 575 ),
( 575 ),
( 575 ),
( 574 ),
( 574 ),
( 574 ),
( 573 ),
( 573 ),
( 573 ),
( 572 ),
( 572 ),
( 572 ),
( 571 ),
( 571 ),
( 571 ),
( 570 ),
( 570 ),
( 570 ),
( 569 ),
( 569 ),
( 569 ),
( 568 ),
( 568 ),
( 567 ),
( 567 ),
( 567 ),
( 566 ),
( 566 ),
( 566 ),
( 565 ),
( 565 ),
( 565 ),
( 564 ),
( 564 ),
( 564 ),
( 563 ),
( 563 ),
( 563 ),
( 562 ),
( 562 ),
( 562 ),
( 561 ),
( 561 ),
( 561 ),
( 560 ),
( 560 ),
( 560 ),
( 559 ),
( 559 ),
( 559 ),
( 558 ),
( 558 ),
( 558 ),
( 557 ),
( 557 ),
( 557 ),
( 556 ),
( 556 ),
( 556 ),
( 555 ),
( 555 ),
( 555 ),
( 554 ),
( 554 ),
( 554 ),
( 553 ),
( 553 ),
( 553 ),
( 552 ),
( 552 ),
( 551 ),
( 551 ),
( 551 ),
( 550 ),
( 550 ),
( 550 ),
( 549 ),
( 549 ),
( 549 ),
( 548 ),
( 548 ),
( 548 ),
( 547 ),
( 547 ),
( 547 ),
( 546 ),
( 546 ),
( 546 ),
( 545 ),
( 545 ),
( 545 ),
( 544 ),
( 544 ),
( 544 ),
( 543 ),
( 543 ),
( 543 ),
( 542 ),
( 542 ),
( 542 ),
( 541 ),
( 541 ),
( 541 ),
( 540 ),
( 540 ),
( 540 ),
( 539 ),
( 539 ),
( 539 ),
( 538 ),
( 538 ),
( 538 ),
( 537 ),
( 537 ),
( 536 ),
( 536 ),
( 536 ),
( 535 ),
( 535 ),
( 535 ),
( 534 ),
( 534 ),
( 534 ),
( 533 ),
( 533 ),
( 533 ),
( 532 ),
( 532 ),
( 532 ),
( 531 ),
( 531 ),
( 531 ),
( 530 ),
( 530 ),
( 530 ),
( 529 ),
( 529 ),
( 529 ),
( 528 ),
( 528 ),
( 528 ),
( 527 ),
( 527 ),
( 527 ),
( 526 ),
( 526 ),
( 526 ),
( 525 ),
( 525 ),
( 525 ),
( 524 ),
( 524 ),
( 524 ),
( 523 ),
( 523 ),
( 523 ),
( 522 ),
( 522 ),
( 522 ),
( 521 ),
( 521 ),
( 521 ),
( 520 ),
( 520 ),
( 520 ),
( 519 ),
( 519 ),
( 519 ),
( 518 ),
( 518 ),
( 518 ),
( 517 ),
( 517 ),
( 516 ),
( 516 ),
( 516 ),
( 515 ),
( 515 ),
( 515 ),
( 514 ),
( 514 ),
( 514 ),
( 513 ),
( 513 ),
( 513 ),
( 512 ),
( 512 ),
( 512 ),
( 511 ),
( 511 ),
( 511 ),
( 510 ),
( 510 ),
( 510 ),
( 509 ),
( 509 ),
( 509 ),
( 508 ),
( 508 ),
( 508 ),
( 508 ),
( 507 ),
( 507 ),
( 507 ),
( 506 ),
( 506 ),
( 506 ),
( 505 ),
( 505 ),
( 505 ),
( 504 ),
( 504 ),
( 504 ),
( 503 ),
( 503 ),
( 503 ),
( 502 ),
( 502 ),
( 502 ),
( 501 ),
( 501 ),
( 501 ),
( 500 ),
( 500 ),
( 500 ),
( 499 ),
( 499 ),
( 499 ),
( 498 ),
( 498 ),
( 498 ),
( 497 ),
( 497 ),
( 497 ),
( 496 ),
( 496 ),
( 496 ),
( 495 ),
( 495 ),
( 495 ),
( 494 ),
( 494 ),
( 494 ),
( 494 ),
( 493 ),
( 493 ),
( 493 ),
( 492 ),
( 492 ),
( 492 ),
( 491 ),
( 491 ),
( 491 ),
( 490 ),
( 490 ),
( 490 ),
( 489 ),
( 489 ),
( 489 ),
( 488 ),
( 488 ),
( 488 ),
( 487 ),
( 487 ),
( 487 ),
( 487 ),
( 486 ),
( 486 ),
( 486 ),
( 485 ),
( 485 ),
( 485 ),
( 484 ),
( 484 ),
( 484 ),
( 483 ),
( 483 ),
( 483 ),
( 483 ),
( 482 ),
( 482 ),
( 482 ),
( 481 ),
( 481 ),
( 481 ),
( 480 ),
( 480 ),
( 480 ),
( 479 ),
( 479 ),
( 479 ),
( 479 ),
( 478 ),
( 478 ),
( 478 ),
( 477 ),
( 477 ),
( 477 ),
( 476 ),
( 476 ),
( 476 ),
( 476 ),
( 475 ),
( 475 ),
( 475 ),
( 474 ),
( 474 ),
( 474 ),
( 473 ),
( 473 ),
( 473 ),
( 473 ),
( 472 ),
( 472 ),
( 472 ),
( 471 ),
( 471 ),
( 471 ),
( 471 ),
( 470 ),
( 470 ),
( 470 ),
( 469 ),
( 469 ),
( 469 ),
( 469 ),
( 468 ),
( 468 ),
( 468 ),
( 467 ),
( 467 ),
( 467 ),
( 467 ),
( 466 ),
( 466 ),
( 466 ),
( 465 ),
( 465 ),
( 465 ),
( 465 ),
( 464 ),
( 464 ),
( 464 ),
( 463 ),
( 463 ),
( 463 ),
( 463 ),
( 462 ),
( 462 ),
( 462 ),
( 461 ),
( 461 ),
( 461 ),
( 461 ),
( 460 ),
( 460 ),
( 460 ),
( 460 ),
( 459 ),
( 459 ),
( 459 ),
( 458 ),
( 458 ),
( 458 ),
( 458 ),
( 457 ),
( 457 ),
( 457 ),
( 457 ),
( 456 ),
( 456 ),
( 456 ),
( 456 ),
( 455 ),
( 455 ),
( 455 ),
( 455 ),
( 454 ),
( 454 ),
( 454 ),
( 453 ),
( 453 ),
( 453 ),
( 453 ),
( 452 ),
( 452 ),
( 452 ),
( 452 ),
( 451 ),
( 451 ),
( 451 ),
( 451 ),
( 450 ),
( 450 ),
( 450 ),
( 450 ),
( 449 ),
( 449 ),
( 449 ),
( 449 ),
( 448 ),
( 448 ),
( 448 ),
( 448 ),
( 447 ),
( 447 ),
( 447 ),
( 447 ),
( 447 ),
( 446 ),
( 446 ),
( 446 ),
( 446 ),
( 445 ),
( 445 ),
( 445 ),
( 445 ),
( 444 ),
( 444 ),
( 444 ),
( 444 ),
( 443 ),
( 443 ),
( 443 ),
( 443 ),
( 442 ),
( 442 ),
( 442 ),
( 442 ),
( 442 ),
( 441 ),
( 441 ),
( 441 ),
( 441 ),
( 440 ),
( 440 ),
( 440 ),
( 440 ),
( 440 ),
( 439 ),
( 439 ),
( 439 ),
( 439 ),
( 438 ),
( 438 ),
( 438 ),
( 438 ),
( 438 ),
( 437 ),
( 437 ),
( 437 ),
( 437 ),
( 436 ),
( 436 ),
( 436 ),
( 436 ),
( 436 ),
( 435 ),
( 435 ),
( 435 ),
( 435 ),
( 435 ),
( 434 ),
( 434 ),
( 434 ),
( 434 ),
( 434 ),
( 433 ),
( 433 ),
( 433 ),
( 433 ),
( 433 ),
( 432 ),
( 432 ),
( 432 ),
( 432 ),
( 432 ),
( 431 ),
( 431 ),
( 431 ),
( 431 ),
( 431 ),
( 430 ),
( 430 ),
( 430 ),
( 430 ),
( 430 ),
( 429 ),
( 429 ),
( 429 ),
( 429 ),
( 429 ),
( 428 ),
( 428 ),
( 428 ),
( 428 ),
( 428 ),
( 427 ),
( 427 ),
( 427 ),
( 427 ),
( 427 ),
( 427 ),
( 426 ),
( 426 ),
( 426 ),
( 426 ),
( 426 ),
( 425 ),
( 425 ),
( 425 ),
( 425 ),
( 425 ),
( 425 ),
( 424 ),
( 424 ),
( 424 ),
( 424 ),
( 424 ),
( 424 ),
( 423 ),
( 423 ),
( 423 ),
( 423 ),
( 423 ),
( 422 ),
( 422 ),
( 422 ),
( 422 ),
( 422 ),
( 422 ),
( 421 ),
( 421 ),
( 421 ),
( 421 ),
( 421 ),
( 421 ),
( 420 ),
( 420 ),
( 420 ),
( 420 ),
( 420 ),
( 420 ),
( 419 ),
( 419 ),
( 419 ),
( 419 ),
( 419 ),
( 419 ),
( 419 ),
( 418 ),
( 418 ),
( 418 ),
( 418 ),
( 418 ),
( 418 ),
( 417 ),
( 417 ),
( 417 ),
( 417 ),
( 417 ),
( 417 ),
( 416 ),
( 416 ),
( 416 ),
( 416 ),
( 416 ),
( 416 ),
( 416 ),
( 415 ),
( 415 ),
( 415 ),
( 415 ),
( 415 ),
( 415 ),
( 415 ),
( 414 ),
( 414 ),
( 414 ),
( 414 ),
( 414 ),
( 414 ),
( 413 ),
( 413 ),
( 413 ),
( 413 ),
( 413 ),
( 413 ),
( 413 ),
( 412 ),
( 412 ),
( 412 ),
( 412 ),
( 412 ),
( 412 ),
( 412 ),
( 411 ),
( 411 ),
( 411 ),
( 411 ),
( 411 ),
( 411 ),
( 411 ),
( 410 ),
( 410 ),
( 410 ),
( 410 ),
( 410 ),
( 410 ),
( 410 ),
( 409 ),
( 409 ),
( 409 ),
( 409 ),
( 409 ),
( 409 ),
( 409 ),
( 408 ),
( 408 ),
( 408 ),
( 408 ),
( 408 ),
( 408 ),
( 408 ),
( 407 ),
( 407 ),
( 407 ),
( 407 ),
( 407 ),
( 407 ),
( 407 ),
( 406 ),
( 406 ),
( 406 ),
( 406 ),
( 406 ),
( 406 ),
( 405 ),
( 405 ),
( 405 ),
( 405 ),
( 405 ),
( 405 ),
( 405 ),
( 404 ),
( 404 ),
( 404 ),
( 404 ),
( 404 ),
( 404 ),
( 404 ),
( 403 ),
( 403 ),
( 403 ),
( 403 ),
( 403 ),
( 403 ),
( 403 ),
( 402 ),
( 402 ),
( 402 ),
( 402 ),
( 402 ),
( 402 ),
( 401 ),
( 401 ),
( 401 ),
( 401 ),
( 401 ),
( 401 ),
( 401 ),
( 400 ),
( 400 ),
( 400 ),
( 400 ),
( 400 ),
( 400 ),
( 399 ),
( 399 ),
( 399 ),
( 399 ),
( 399 ),
( 399 ),
( 398 ),
( 398 ),
( 398 ),
( 398 ),
( 398 ),
( 398 ),
( 397 ),
( 397 ),
( 397 ),
( 397 ),
( 397 ),
( 397 ),
( 396 ),
( 396 ),
( 396 ),
( 396 ),
( 396 ),
( 395 ),
( 395 ),
( 395 ),
( 395 ),
( 395 ),
( 395 ),
( 394 ),
( 394 ),
( 394 ),
( 394 ),
( 394 ),
( 393 ),
( 393 ),
( 393 ),
( 393 ),
( 393 ),
( 392 ),
( 392 ),
( 392 ),
( 392 ),
( 392 ),
( 391 ),
( 391 ),
( 391 ),
( 391 ),
( 391 ),
( 390 ),
( 390 ),
( 390 ),
( 390 ),
( 390 ),
( 389 ),
( 389 ),
( 389 ),
( 389 ),
( 388 ),
( 388 ),
( 388 ),
( 388 ),
( 388 ),
( 387 ),
( 387 ),
( 387 ),
( 387 ),
( 386 ),
( 386 ),
( 386 ),
( 386 ),
( 385 ),
( 385 ),
( 385 ),
( 385 ),
( 384 ),
( 384 ),
( 384 ),
( 384 ),
( 383 ),
( 383 ),
( 383 ),
( 383 ),
( 382 ),
( 382 ),
( 382 ),
( 381 ),
( 381 ),
( 381 ),
( 381 ),
( 380 ),
( 380 ),
( 380 ),
( 379 ),
( 379 ),
( 379 ),
( 379 ),
( 378 ),
( 378 ),
( 378 ),
( 377 ),
( 377 ),
( 377 ),
( 376 ),
( 376 ),
( 376 ),
( 375 ),
( 375 ),
( 375 ),
( 374 ),
( 374 ),
( 374 ),
( 373 ),
( 373 ),
( 373 ),
( 372 ),
( 372 ),
( 372 ),
( 371 ),
( 371 ),
( 371 ),
( 370 ),
( 370 ),
( 369 ),
( 369 ),
( 369 ),
( 368 ),
( 368 ),
( 367 ),
( 367 ),
( 367 ),
( 366 ),
( 366 ),
( 365 ),
( 365 ),
( 365 ),
( 364 ),
( 364 ),
( 363 ),
( 363 ),
( 363 ),
( 362 ),
( 362 ),
( 361 ),
( 361 ),
( 360 ),
( 360 ),
( 359 ),
( 359 ),
( 358 ),
( 358 ),
( 358 ),
( 357 ),
( 357 ),
( 356 ),
( 356 ),
( 355 ),
( 355 ),
( 354 ),
( 354 ),
( 353 ),
( 353 ),
( 352 ),
( 352 ),
( 351 ),
( 350 ),
( 350 ),
( 349 ),
( 349 ),
( 348 ),
( 348 ),
( 347 ),
( 347 ),
( 346 ),
( 345 ),
( 345 ),
( 344 ),
( 344 ),
( 343 ),
( 342 ),
( 342 ),
( 341 ),
( 341 ),
( 340 ),
( 339 ),
( 339 ),
( 338 ),
( 338 ),
( 337 ),
( 336 ),
( 336 ),
( 335 ),
( 334 ),
( 334 ),
( 333 ),
( 332 ),
( 332 ),
( 331 ),
( 330 ),
( 329 ),
( 329 ),
( 328 ),
( 327 ),
( 327 ),
( 326 ),
( 325 ),
( 324 ),
( 324 ),
( 323 ),
( 322 ),
( 321 ),
( 320 ),
( 320 ),
( 319 ),
( 318 ),
( 317 ),
( 316 ),
( 316 ),
( 315 ),
( 314 ),
( 313 ),
( 312 ),
( 311 ),
( 311 ),
( 310 ),
( 309 ),
( 308 ),
( 307 ),
( 306 ),
( 305 ),
( 304 ),
( 304 ),
( 303 ),
( 302 ),
( 301 ),
( 300 ),
( 299 ),
( 298 ),
( 297 ),
( 296 ),
( 295 ),
( 294 ),
( 293 ),
( 292 ),
( 291 ),
( 290 ),
( 289 ),
( 288 ),
( 287 ),
( 286 ),
( 285 ),
( 284 ),
( 283 ),
( 282 ),
( 281 ),
( 279 ),
( 278 ),
( 277 ),
( 276 ),
( 275 ),
( 274 ),
( 273 ),
( 272 ),
( 270 ),
( 269 ),
( 268 ),
( 267 ),
( 266 ),
( 264 ),
( 263 ),
( 262 ),
( 261 ),
( 259 ),
( 258 ),
( 257 ),
( 256 ),
( 254 ),
( 253 ),
( 252 ),
( 251 ),
( 249 ),
( 248 ),
( 247 ),
( 245 ),
( 244 ),
( 242 ),
( 241 ),
( 240 ),
( 238 ),
( 237 ),
( 235 ),
( 234 ),
( 233 ),
( 231 ),
( 230 ),
( 228 ),
( 227 ),
( 225 ),
( 224 ),
( 222 ),
( 221 ),
( 219 ),
( 218 ),
( 216 ),
( 214 ),
( 213 ),
( 211 ),
( 210 ),
( 208 ),
( 206 ),
( 205 ),
( 203 ),
( 201 ),
( 200 ),
( 198 ),
( 196 ),
( 195 ),
( 193 ),
( 191 ),
( 190 ),
( 188 ),
( 186 ),
( 184 ),
( 182 ),
( 181 ),
( 179 ),
( 177 ),
( 175 ),
( 173 ),
( 171 ),
( 170 ),
( 168 ),
( 166 ),
( 164 ),
( 162 ),
( 160 ),
( 158 ),
( 156 ),
( 154 ),
( 152 ),
( 150 ),
( 148 ),
( 146 ),
( 144 ),
( 142 ),
( 140 ),
( 138 ),
( 136 ),
( 133 ),
( 131 ),
( 129 ),
( 127 ),
( 125 ),
( 123 ),
( 120 ),
( 118 ),
( 116 ),
( 114 ),
( 111 ),
( 109 ),
( 107 ),
( 104 ),
( 102 ),
( 100 ),
( 97 ),
( 95 ),
( 93 ),
( 90 ),
( 88 ),
( 85 ),
( 83 ),
( 80 ),
( 78 ),
( 75 ),
( 73 ),
( 70 ),
( 68 ),
( 65 ),
( 63 ),
( 60 ),
( 58 ),
( 55 ),
( 52 ),
( 50 ),
( 47 ),
( 44 ),
( 41 ),
( 39 ),
( 36 ),
( 33 ),
( 30 ),
( 28 ),
( 25 ),
( 22 ),
( 19 ),
( 16 ),
( 13 ),
( 10 ),
( 7 ),
( 5 ),
( 2 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 ),
( 0 )





);


begin    	

   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));

end behavior;
